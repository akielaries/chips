module alu_4_bit
